module deco ( 
	clr,
	clk,
	u,
	d,
	display,
	contanillo
	) ;

input  clr;
input  clk;
input [3:0] u;
input [2:0] d;
inout [6:0] display;
inout [2:0] contanillo;
