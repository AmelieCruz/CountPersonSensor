module detector ( 
	clr,
	clk,
	sen,
	d,
	u
	) ;

input  clr;
input  clk;
input [1:0] sen;
inout [2:0] d;
inout [3:0] u;
